/* 
Guia_0804.v 
855842 - Mateus Resende Ottoni

iverilog -o Guia_0804.vvp Guia_0804.v
vvp Guia_0804.vvp
*/



// Desigualdade
//----------------------------------------
module inequal (output s,
                   input a, b, c);

// Dados locais
wire w1;

// Processo
xor	XOR  (  w1,   a,   b);
or	OR   (   s,  w1,   c); // Saída


endmodule
//----------------------------------------

// Modulo de desigualdade
//----------------------------------------
module f04 (output s,
            input  a0, b0, a1, b1,
                   a2, b2, a3, b3);

// Dados locais
reg valor0 = 1'b0;
wire res01, res02, res03;

// Processo
inequal IN1 ( res01, a0, b0, valor0);
inequal IN2 ( res02, a1, b1,  res01);
inequal IN3 ( res03, a2, b2,  res02);
inequal IN4 (     s, a3, b3,  res03); // Saída

endmodule
//----------------------------------------




// Modulo principal
module Guia_0804; 

// Definir dados
reg a0, b0, a1, b1, a2, b2, a3, b3;
wire w;

f04    f04_ ( w,
              a0, b0, a1, b1, a2, b2, a3, b3);


 initial
  begin
   a0     = 1'b0;
   b0     = 1'b0;
   a1     = 1'b0;
   b1     = 1'b0;
   a2     = 1'b0;
   b2     = 1'b0;
   a3     = 1'b0;
   b3     = 1'b0;
  end


// Main 
initial 
begin : main 

$display ( "Guia_0804" );

/*	Mostrar valores em tabela				*/
$display ( "" );
$display ( "_________________________________" );
$display ( "||    a |    b || desigualdade ||" );
$display ( "||------|------||--------------||" );
$monitor ( "|| %b%b%b%b | %b%b%b%b ||            %b ||",
              a3, a2, a1, a0,
                         b3, b2, b1, b0,
                                                  w );
/*								*/

/*	Atualizar valores ( a = 00)	*/

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 01)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 02)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 03)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 04)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 05)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 06)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 07)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 08)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b0; a3 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 09)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 10)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 11)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 12)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 13)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 14)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 15)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/



end // main 

endmodule // Guia_0804

/*	Previsão de Testes 		*/
/*


_________________________________
||    a |    b || desigualdade ||
||------|------||--------------||
|| 0000 | 0000 ||            0 ||
|| 0000 | 0001 ||            1 ||
|| 0000 | 0010 ||            1 ||
|| 0000 | 0011 ||            1 ||
|| 0000 | 0100 ||            1 ||
|| 0000 | 0101 ||            1 ||
|| 0000 | 0110 ||            1 ||
|| 0000 | 0111 ||            1 ||
|| 0000 | 1000 ||            1 ||
|| 0000 | 1001 ||            1 ||
|| 0000 | 1010 ||            1 ||
|| 0000 | 1011 ||            1 ||
|| 0000 | 1100 ||            1 ||
|| 0000 | 1101 ||            1 ||
|| 0000 | 1110 ||            1 ||
|| 0000 | 1111 ||            1 ||
|| 0001 | 0000 ||            1 ||
|| 0001 | 0001 ||            0 ||
|| 0001 | 0010 ||            1 ||
|| 0001 | 0011 ||            1 ||
|| 0001 | 0100 ||            1 ||
|| 0001 | 0101 ||            1 ||
|| 0001 | 0110 ||            1 ||
|| 0001 | 0111 ||            1 ||
|| 0001 | 1000 ||            1 ||
|| 0001 | 1001 ||            1 ||
|| 0001 | 1010 ||            1 ||
|| 0001 | 1011 ||            1 ||
|| 0001 | 1100 ||            1 ||
|| 0001 | 1101 ||            1 ||
|| 0001 | 1110 ||            1 ||
|| 0001 | 1111 ||            1 ||
|| 0010 | 0000 ||            1 ||
|| 0010 | 0001 ||            1 ||
|| 0010 | 0010 ||            0 ||
|| 0010 | 0011 ||            1 ||
|| 0010 | 0100 ||            1 ||
|| 0010 | 0101 ||            1 ||
|| 0010 | 0110 ||            1 ||
|| 0010 | 0111 ||            1 ||
|| 0010 | 1000 ||            1 ||
|| 0010 | 1001 ||            1 ||
|| 0010 | 1010 ||            1 ||
|| 0010 | 1011 ||            1 ||
|| 0010 | 1100 ||            1 ||
|| 0010 | 1101 ||            1 ||
|| 0010 | 1110 ||            1 ||
|| 0010 | 1111 ||            1 ||
|| 0011 | 0000 ||            1 ||
|| 0011 | 0001 ||            1 ||
|| 0011 | 0010 ||            1 ||
|| 0011 | 0011 ||            0 ||
|| 0011 | 0100 ||            1 ||
|| 0011 | 0101 ||            1 ||
|| 0011 | 0110 ||            1 ||
|| 0011 | 0111 ||            1 ||
|| 0011 | 1000 ||            1 ||
|| 0011 | 1001 ||            1 ||
|| 0011 | 1010 ||            1 ||
|| 0011 | 1011 ||            1 ||
|| 0011 | 1100 ||            1 ||
|| 0011 | 1101 ||            1 ||
|| 0011 | 1110 ||            1 ||
|| 0011 | 1111 ||            1 ||
|| 0100 | 0000 ||            1 ||
|| 0100 | 0001 ||            1 ||
|| 0100 | 0010 ||            1 ||
|| 0100 | 0011 ||            1 ||
|| 0100 | 0100 ||            0 ||
|| 0100 | 0101 ||            1 ||
|| 0100 | 0110 ||            1 ||
|| 0100 | 0111 ||            1 ||
|| 0100 | 1000 ||            1 ||
|| 0100 | 1001 ||            1 ||
|| 0100 | 1010 ||            1 ||
|| 0100 | 1011 ||            1 ||
|| 0100 | 1100 ||            1 ||
|| 0100 | 1101 ||            1 ||
|| 0100 | 1110 ||            1 ||
|| 0100 | 1111 ||            1 ||
|| 0101 | 0000 ||            1 ||
|| 0101 | 0001 ||            1 ||
|| 0101 | 0010 ||            1 ||
|| 0101 | 0011 ||            1 ||
|| 0101 | 0100 ||            1 ||
|| 0101 | 0101 ||            0 ||
|| 0101 | 0110 ||            1 ||
|| 0101 | 0111 ||            1 ||
|| 0101 | 1000 ||            1 ||
|| 0101 | 1001 ||            1 ||
|| 0101 | 1010 ||            1 ||
|| 0101 | 1011 ||            1 ||
|| 0101 | 1100 ||            1 ||
|| 0101 | 1101 ||            1 ||
|| 0101 | 1110 ||            1 ||
|| 0101 | 1111 ||            1 ||
|| 0110 | 0000 ||            1 ||
|| 0110 | 0001 ||            1 ||
|| 0110 | 0010 ||            1 ||
|| 0110 | 0011 ||            1 ||
|| 0110 | 0100 ||            1 ||
|| 0110 | 0101 ||            1 ||
|| 0110 | 0110 ||            0 ||
|| 0110 | 0111 ||            1 ||
|| 0110 | 1000 ||            1 ||
|| 0110 | 1001 ||            1 ||
|| 0110 | 1010 ||            1 ||
|| 0110 | 1011 ||            1 ||
|| 0110 | 1100 ||            1 ||
|| 0110 | 1101 ||            1 ||
|| 0110 | 1110 ||            1 ||
|| 0110 | 1111 ||            1 ||
|| 0111 | 0000 ||            1 ||
|| 0111 | 0001 ||            1 ||
|| 0111 | 0010 ||            1 ||
|| 0111 | 0011 ||            1 ||
|| 0111 | 0100 ||            1 ||
|| 0111 | 0101 ||            1 ||
|| 0111 | 0110 ||            1 ||
|| 0111 | 0111 ||            0 ||
|| 0111 | 1000 ||            1 ||
|| 0111 | 1001 ||            1 ||
|| 0111 | 1010 ||            1 ||
|| 0111 | 1011 ||            1 ||
|| 0111 | 1100 ||            1 ||
|| 0111 | 1101 ||            1 ||
|| 0111 | 1110 ||            1 ||
|| 0111 | 1111 ||            1 ||
|| 1000 | 0000 ||            1 ||
|| 1000 | 0001 ||            1 ||
|| 1000 | 0010 ||            1 ||
|| 1000 | 0011 ||            1 ||
|| 1000 | 0100 ||            1 ||
|| 1000 | 0101 ||            1 ||
|| 1000 | 0110 ||            1 ||
|| 1000 | 0111 ||            1 ||
|| 1000 | 1000 ||            0 ||
|| 1000 | 1001 ||            1 ||
|| 1000 | 1010 ||            1 ||
|| 1000 | 1011 ||            1 ||
|| 1000 | 1100 ||            1 ||
|| 1000 | 1101 ||            1 ||
|| 1000 | 1110 ||            1 ||
|| 1000 | 1111 ||            1 ||
|| 1001 | 0000 ||            1 ||
|| 1001 | 0001 ||            1 ||
|| 1001 | 0010 ||            1 ||
|| 1001 | 0011 ||            1 ||
|| 1001 | 0100 ||            1 ||
|| 1001 | 0101 ||            1 ||
|| 1001 | 0110 ||            1 ||
|| 1001 | 0111 ||            1 ||
|| 1001 | 1000 ||            1 ||
|| 1001 | 1001 ||            0 ||
|| 1001 | 1010 ||            1 ||
|| 1001 | 1011 ||            1 ||
|| 1001 | 1100 ||            1 ||
|| 1001 | 1101 ||            1 ||
|| 1001 | 1110 ||            1 ||
|| 1001 | 1111 ||            1 ||
|| 1010 | 0000 ||            1 ||
|| 1010 | 0001 ||            1 ||
|| 1010 | 0010 ||            1 ||
|| 1010 | 0011 ||            1 ||
|| 1010 | 0100 ||            1 ||
|| 1010 | 0101 ||            1 ||
|| 1010 | 0110 ||            1 ||
|| 1010 | 0111 ||            1 ||
|| 1010 | 1000 ||            1 ||
|| 1010 | 1001 ||            1 ||
|| 1010 | 1010 ||            0 ||
|| 1010 | 1011 ||            1 ||
|| 1010 | 1100 ||            1 ||
|| 1010 | 1101 ||            1 ||
|| 1010 | 1110 ||            1 ||
|| 1010 | 1111 ||            1 ||
|| 1011 | 0000 ||            1 ||
|| 1011 | 0001 ||            1 ||
|| 1011 | 0010 ||            1 ||
|| 1011 | 0011 ||            1 ||
|| 1011 | 0100 ||            1 ||
|| 1011 | 0101 ||            1 ||
|| 1011 | 0110 ||            1 ||
|| 1011 | 0111 ||            1 ||
|| 1011 | 1000 ||            1 ||
|| 1011 | 1001 ||            1 ||
|| 1011 | 1010 ||            1 ||
|| 1011 | 1011 ||            0 ||
|| 1011 | 1100 ||            1 ||
|| 1011 | 1101 ||            1 ||
|| 1011 | 1110 ||            1 ||
|| 1011 | 1111 ||            1 ||
|| 1100 | 0000 ||            1 ||
|| 1100 | 0001 ||            1 ||
|| 1100 | 0010 ||            1 ||
|| 1100 | 0011 ||            1 ||
|| 1100 | 0100 ||            1 ||
|| 1100 | 0101 ||            1 ||
|| 1100 | 0110 ||            1 ||
|| 1100 | 0111 ||            1 ||
|| 1100 | 1000 ||            1 ||
|| 1100 | 1001 ||            1 ||
|| 1100 | 1010 ||            1 ||
|| 1100 | 1011 ||            1 ||
|| 1100 | 1100 ||            0 ||
|| 1100 | 1101 ||            1 ||
|| 1100 | 1110 ||            1 ||
|| 1100 | 1111 ||            1 ||
|| 1101 | 0000 ||            1 ||
|| 1101 | 0001 ||            1 ||
|| 1101 | 0010 ||            1 ||
|| 1101 | 0011 ||            1 ||
|| 1101 | 0100 ||            1 ||
|| 1101 | 0101 ||            1 ||
|| 1101 | 0110 ||            1 ||
|| 1101 | 0111 ||            1 ||
|| 1101 | 1000 ||            1 ||
|| 1101 | 1001 ||            1 ||
|| 1101 | 1010 ||            1 ||
|| 1101 | 1011 ||            1 ||
|| 1101 | 1100 ||            1 ||
|| 1101 | 1101 ||            0 ||
|| 1101 | 1110 ||            1 ||
|| 1101 | 1111 ||            1 ||
|| 1110 | 0000 ||            1 ||
|| 1110 | 0001 ||            1 ||
|| 1110 | 0010 ||            1 ||
|| 1110 | 0011 ||            1 ||
|| 1110 | 0100 ||            1 ||
|| 1110 | 0101 ||            1 ||
|| 1110 | 0110 ||            1 ||
|| 1110 | 0111 ||            1 ||
|| 1110 | 1000 ||            1 ||
|| 1110 | 1001 ||            1 ||
|| 1110 | 1010 ||            1 ||
|| 1110 | 1011 ||            1 ||
|| 1110 | 1100 ||            1 ||
|| 1110 | 1101 ||            1 ||
|| 1110 | 1110 ||            0 ||
|| 1110 | 1111 ||            1 ||
|| 1111 | 0000 ||            1 ||
|| 1111 | 0001 ||            1 ||
|| 1111 | 0010 ||            1 ||
|| 1111 | 0011 ||            1 ||
|| 1111 | 0100 ||            1 ||
|| 1111 | 0101 ||            1 ||
|| 1111 | 0110 ||            1 ||
|| 1111 | 0111 ||            1 ||
|| 1111 | 1000 ||            1 ||
|| 1111 | 1001 ||            1 ||
|| 1111 | 1010 ||            1 ||
|| 1111 | 1011 ||            1 ||
|| 1111 | 1100 ||            1 ||
|| 1111 | 1101 ||            1 ||
|| 1111 | 1110 ||            1 ||
|| 1111 | 1111 ||            0 ||


*/
/*					*/
