/* 
Guia_0801.v 
855842 - Mateus Resende Ottoni

iverilog -o Guia_0801.vvp Guia_0801.v
vvp Guia_0801.vvp
*/



// Meia Soma
//----------------------------------------
module half_adder (output s0, output s1,
                   input a, b);

// Saída 1
   xor XOR (	s0,	a,	b);

// Saída 2
   and AND (	s1,	a,	b);

endmodule
//----------------------------------------

// Soma completa
//----------------------------------------
module full_adder (output s0, output s1,
                   input a, b, c);

// Dados locais
wire w01, w11, w12;

// Processo
half_adder HA1 ( w01, w11,   a,   b);
half_adder HA2 (  s1, w12, w01,   c); // Saída s1
or         OR  (  s0,      w11, w12); // Saída s0



endmodule
//----------------------------------------

// Modulo de soma
//----------------------------------------
module f01 (output s1, output s2, output s3,
            output s4, output s5,
            input  a0, b0, a1, b1,
                   a2, b2, a3, b3);

// Dados locais
reg valor0 = 1'b0;
wire res01, res02, res03;

// Processo
full_adder FA1 ( res01, s1, a0, b0, valor0); // Saída s1
full_adder FA2 ( res02, s2, a1, b1,  res01); // Saída s2
full_adder FA3 ( res03, s3, a2, b2,  res02); // Saída s3
full_adder FA4 (    s5, s4, a3, b3,  res03); // Saída s4 e s5

endmodule
//----------------------------------------




// Modulo principal
module Guia_0801; 

// Definir dados
reg a0, b0, a1, b1, a2, b2, a3, b3;
wire w1, w2, w3, w4, w5;

f01    f01_ (w1, w2, w3, w4, w5,
             a0, b0, a1, b1, a2, b2, a3, b3);


 initial
  begin
   a0     = 1'b0;
   b0     = 1'b0;
   a1     = 1'b0;
   b1     = 1'b0;
   a2     = 1'b0;
   b2     = 1'b0;
   a3     = 1'b0;
   b3     = 1'b0;
  end


// Main 
initial 
begin : main 

$display ( "Guia_0801" );

/*	Mostrar valores em tabela				*/
$display ( "" );
$display ( "______________________________" );
$display ( "||    a |    b ||   soma   ||" );
$display ( "||------|------||----------||" );
$monitor ( "|| %b%b%b%b | %b%b%b%b ||    %b%b%b%b%b ||",
              a3, a2, a1, a0,
                         b3, b2, b1, b0,
                                     w5, w4, w3, w2, w1 );
/*								*/

/*	Atualizar valores ( a = 00)	*/

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 01)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 02)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 03)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 04)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 05)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 06)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 07)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 08)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b0; a3 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 09)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 10)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 11)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 12)	*/

#1;  a0 = 1'b0; a1 = 1'b0; a2 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 13)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 14)	*/

#1;  a0 = 1'b0; a1 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/

/*	Atualizar valores ( a = 15)	*/

#1;  a0 = 1'b1;
     b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b0;

#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b0; b3 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b0; b2 = 1'b1;
#1;  b0 = 1'b1;
#1;  b0 = 1'b0; b1 = 1'b1;
#1;  b0 = 1'b1;

/*					*/



end // main 

endmodule // Guia_0801

/*	Previsão de Testes 		*/
/*


______________________________
||    a |    b || resultado ||
||------|------||-----------||
|| 0000 | 0000 ||     00000 ||
|| 0000 | 0001 ||     00001 ||
|| 0000 | 0010 ||     00010 ||
|| 0000 | 0011 ||     00011 ||
|| 0000 | 0100 ||     00100 ||
|| 0000 | 0101 ||     00101 ||
|| 0000 | 0110 ||     00110 ||
|| 0000 | 0111 ||     00111 ||
|| 0000 | 1000 ||     01000 ||
|| 0000 | 1001 ||     01001 ||
|| 0000 | 1010 ||     01010 ||
|| 0000 | 1011 ||     01011 ||
|| 0000 | 1100 ||     01100 ||
|| 0000 | 1101 ||     01101 ||
|| 0000 | 1110 ||     01110 ||
|| 0000 | 1111 ||     01111 ||
|| 0001 | 0000 ||     00001 ||
|| 0001 | 0001 ||     00010 ||
|| 0001 | 0010 ||     00011 ||
|| 0001 | 0011 ||     00100 ||
|| 0001 | 0100 ||     00101 ||
|| 0001 | 0101 ||     00110 ||
|| 0001 | 0110 ||     00111 ||
|| 0001 | 0111 ||     01000 ||
|| 0001 | 1000 ||     01001 ||
|| 0001 | 1001 ||     01010 ||
|| 0001 | 1010 ||     01011 ||
|| 0001 | 1011 ||     01100 ||
|| 0001 | 1100 ||     01101 ||
|| 0001 | 1101 ||     01110 ||
|| 0001 | 1110 ||     01111 ||
|| 0001 | 1111 ||     10000 ||
|| 0010 | 0000 ||     00010 ||
|| 0010 | 0001 ||     00011 ||
|| 0010 | 0010 ||     00100 ||
|| 0010 | 0011 ||     00101 ||
|| 0010 | 0100 ||     00110 ||
|| 0010 | 0101 ||     00111 ||
|| 0010 | 0110 ||     01000 ||
|| 0010 | 0111 ||     01001 ||
|| 0010 | 1000 ||     01010 ||
|| 0010 | 1001 ||     01011 ||
|| 0010 | 1010 ||     01100 ||
|| 0010 | 1011 ||     01101 ||
|| 0010 | 1100 ||     01110 ||
|| 0010 | 1101 ||     01111 ||
|| 0010 | 1110 ||     10000 ||
|| 0010 | 1111 ||     10001 ||
|| 0011 | 0000 ||     00011 ||
|| 0011 | 0001 ||     00100 ||
|| 0011 | 0010 ||     00101 ||
|| 0011 | 0011 ||     00110 ||
|| 0011 | 0100 ||     00111 ||
|| 0011 | 0101 ||     01000 ||
|| 0011 | 0110 ||     01001 ||
|| 0011 | 0111 ||     01010 ||
|| 0011 | 1000 ||     01011 ||
|| 0011 | 1001 ||     01100 ||
|| 0011 | 1010 ||     01101 ||
|| 0011 | 1011 ||     01110 ||
|| 0011 | 1100 ||     01111 ||
|| 0011 | 1101 ||     10000 ||
|| 0011 | 1110 ||     10001 ||
|| 0011 | 1111 ||     10010 ||
|| 0100 | 0000 ||     00100 ||
|| 0100 | 0001 ||     00101 ||
|| 0100 | 0010 ||     00110 ||
|| 0100 | 0011 ||     00111 ||
|| 0100 | 0100 ||     01000 ||
|| 0100 | 0101 ||     01001 ||
|| 0100 | 0110 ||     01010 ||
|| 0100 | 0111 ||     01011 ||
|| 0100 | 1000 ||     01100 ||
|| 0100 | 1001 ||     01101 ||
|| 0100 | 1010 ||     01110 ||
|| 0100 | 1011 ||     01111 ||
|| 0100 | 1100 ||     10000 ||
|| 0100 | 1101 ||     10001 ||
|| 0100 | 1110 ||     10010 ||
|| 0100 | 1111 ||     10011 ||
|| 0101 | 0000 ||     00101 ||
|| 0101 | 0001 ||     00110 ||
|| 0101 | 0010 ||     00111 ||
|| 0101 | 0011 ||     01000 ||
|| 0101 | 0100 ||     01001 ||
|| 0101 | 0101 ||     01010 ||
|| 0101 | 0110 ||     01011 ||
|| 0101 | 0111 ||     01100 ||
|| 0101 | 1000 ||     01101 ||
|| 0101 | 1001 ||     01110 ||
|| 0101 | 1010 ||     01111 ||
|| 0101 | 1011 ||     10000 ||
|| 0101 | 1100 ||     10001 ||
|| 0101 | 1101 ||     10010 ||
|| 0101 | 1110 ||     10011 ||
|| 0101 | 1111 ||     10100 ||
|| 0110 | 0000 ||     00110 ||
|| 0110 | 0001 ||     00111 ||
|| 0110 | 0010 ||     01000 ||
|| 0110 | 0011 ||     01001 ||
|| 0110 | 0100 ||     01010 ||
|| 0110 | 0101 ||     01011 ||
|| 0110 | 0110 ||     01100 ||
|| 0110 | 0111 ||     01101 ||
|| 0110 | 1000 ||     01110 ||
|| 0110 | 1001 ||     01111 ||
|| 0110 | 1010 ||     10000 ||
|| 0110 | 1011 ||     10001 ||
|| 0110 | 1100 ||     10010 ||
|| 0110 | 1101 ||     10011 ||
|| 0110 | 1110 ||     10100 ||
|| 0110 | 1111 ||     10101 ||
|| 0111 | 0000 ||     00111 ||
|| 0111 | 0001 ||     01000 ||
|| 0111 | 0010 ||     01001 ||
|| 0111 | 0011 ||     01010 ||
|| 0111 | 0100 ||     01011 ||
|| 0111 | 0101 ||     01100 ||
|| 0111 | 0110 ||     01101 ||
|| 0111 | 0111 ||     01110 ||
|| 0111 | 1000 ||     01111 ||
|| 0111 | 1001 ||     10000 ||
|| 0111 | 1010 ||     10001 ||
|| 0111 | 1011 ||     10010 ||
|| 0111 | 1100 ||     10011 ||
|| 0111 | 1101 ||     10100 ||
|| 0111 | 1110 ||     10101 ||
|| 0111 | 1111 ||     10110 ||
|| 1000 | 0000 ||     01000 ||
|| 1000 | 0001 ||     01001 ||
|| 1000 | 0010 ||     01010 ||
|| 1000 | 0011 ||     01011 ||
|| 1000 | 0100 ||     01100 ||
|| 1000 | 0101 ||     01101 ||
|| 1000 | 0110 ||     01110 ||
|| 1000 | 0111 ||     01111 ||
|| 1000 | 1000 ||     10000 ||
|| 1000 | 1001 ||     10001 ||
|| 1000 | 1010 ||     10010 ||
|| 1000 | 1011 ||     10011 ||
|| 1000 | 1100 ||     10100 ||
|| 1000 | 1101 ||     10101 ||
|| 1000 | 1110 ||     10110 ||
|| 1000 | 1111 ||     10111 ||
|| 1001 | 0000 ||     01001 ||
|| 1001 | 0001 ||     01010 ||
|| 1001 | 0010 ||     01011 ||
|| 1001 | 0011 ||     01100 ||
|| 1001 | 0100 ||     01101 ||
|| 1001 | 0101 ||     01110 ||
|| 1001 | 0110 ||     01111 ||
|| 1001 | 0111 ||     10000 ||
|| 1001 | 1000 ||     10001 ||
|| 1001 | 1001 ||     10010 ||
|| 1001 | 1010 ||     10011 ||
|| 1001 | 1011 ||     10100 ||
|| 1001 | 1100 ||     10101 ||
|| 1001 | 1101 ||     10110 ||
|| 1001 | 1110 ||     10111 ||
|| 1001 | 1111 ||     11000 ||
|| 1010 | 0000 ||     01010 ||
|| 1010 | 0001 ||     01011 ||
|| 1010 | 0010 ||     01100 ||
|| 1010 | 0011 ||     01101 ||
|| 1010 | 0100 ||     01110 ||
|| 1010 | 0101 ||     01111 ||
|| 1010 | 0110 ||     10000 ||
|| 1010 | 0111 ||     10001 ||
|| 1010 | 1000 ||     10010 ||
|| 1010 | 1001 ||     10011 ||
|| 1010 | 1010 ||     10100 ||
|| 1010 | 1011 ||     10101 ||
|| 1010 | 1100 ||     10110 ||
|| 1010 | 1101 ||     10111 ||
|| 1010 | 1110 ||     11000 ||
|| 1010 | 1111 ||     11001 ||
|| 1011 | 0000 ||     01011 ||
|| 1011 | 0001 ||     01100 ||
|| 1011 | 0010 ||     01101 ||
|| 1011 | 0011 ||     01110 ||
|| 1011 | 0100 ||     01111 ||
|| 1011 | 0101 ||     10000 ||
|| 1011 | 0110 ||     10001 ||
|| 1011 | 0111 ||     10010 ||
|| 1011 | 1000 ||     10011 ||
|| 1011 | 1001 ||     10100 ||
|| 1011 | 1010 ||     10101 ||
|| 1011 | 1011 ||     10110 ||
|| 1011 | 1100 ||     10111 ||
|| 1011 | 1101 ||     11000 ||
|| 1011 | 1110 ||     11001 ||
|| 1011 | 1111 ||     11010 ||
|| 1100 | 0000 ||     01100 ||
|| 1100 | 0001 ||     01101 ||
|| 1100 | 0010 ||     01110 ||
|| 1100 | 0011 ||     01111 ||
|| 1100 | 0100 ||     10000 ||
|| 1100 | 0101 ||     10001 ||
|| 1100 | 0110 ||     10010 ||
|| 1100 | 0111 ||     10011 ||
|| 1100 | 1000 ||     10100 ||
|| 1100 | 1001 ||     10101 ||
|| 1100 | 1010 ||     10110 ||
|| 1100 | 1011 ||     10111 ||
|| 1100 | 1100 ||     11000 ||
|| 1100 | 1101 ||     11001 ||
|| 1100 | 1110 ||     11010 ||
|| 1100 | 1111 ||     11011 ||
|| 1101 | 0000 ||     01101 ||
|| 1101 | 0001 ||     01110 ||
|| 1101 | 0010 ||     01111 ||
|| 1101 | 0011 ||     10000 ||
|| 1101 | 0100 ||     10001 ||
|| 1101 | 0101 ||     10010 ||
|| 1101 | 0110 ||     10011 ||
|| 1101 | 0111 ||     10100 ||
|| 1101 | 1000 ||     10101 ||
|| 1101 | 1001 ||     10110 ||
|| 1101 | 1010 ||     10111 ||
|| 1101 | 1011 ||     11000 ||
|| 1101 | 1100 ||     11001 ||
|| 1101 | 1101 ||     11010 ||
|| 1101 | 1110 ||     11011 ||
|| 1101 | 1111 ||     11100 ||
|| 1110 | 0000 ||     01110 ||
|| 1110 | 0001 ||     01111 ||
|| 1110 | 0010 ||     10000 ||
|| 1110 | 0011 ||     10001 ||
|| 1110 | 0100 ||     10010 ||
|| 1110 | 0101 ||     10011 ||
|| 1110 | 0110 ||     10100 ||
|| 1110 | 0111 ||     10101 ||
|| 1110 | 1000 ||     10110 ||
|| 1110 | 1001 ||     10111 ||
|| 1110 | 1010 ||     11000 ||
|| 1110 | 1011 ||     11001 ||
|| 1110 | 1100 ||     11010 ||
|| 1110 | 1101 ||     11011 ||
|| 1110 | 1110 ||     11100 ||
|| 1110 | 1111 ||     11101 ||
|| 1111 | 0000 ||     01111 ||
|| 1111 | 0001 ||     10000 ||
|| 1111 | 0010 ||     10001 ||
|| 1111 | 0011 ||     10010 ||
|| 1111 | 0100 ||     10011 ||
|| 1111 | 0101 ||     10100 ||
|| 1111 | 0110 ||     10101 ||
|| 1111 | 0111 ||     10110 ||
|| 1111 | 1000 ||     10111 ||
|| 1111 | 1001 ||     11000 ||
|| 1111 | 1010 ||     11001 ||
|| 1111 | 1011 ||     11010 ||
|| 1111 | 1100 ||     11011 ||
|| 1111 | 1101 ||     11100 ||
|| 1111 | 1110 ||     11101 ||
|| 1111 | 1111 ||     11110 ||


*/
/*					*/
